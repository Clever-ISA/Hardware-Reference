library types;
use types.all;


package alu is

    procedure add_and_scale64(base : in u64, carryin : in u1, index : in u64, scale: in u3, variable carryout : out u1, variable result : out u64) 
    is 
    begin 

    end add_and_scale64;

end alu;