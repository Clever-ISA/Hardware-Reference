library types;
use types.all;

library ieee;
use ieee.std_logic;

architecture clever is
    shared signal clk: std_logic;
end clever;